
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'had2a3c00;
    ram_cell[       1] = 32'h0;  // 32'h43258ffb;
    ram_cell[       2] = 32'h0;  // 32'hfcca45bb;
    ram_cell[       3] = 32'h0;  // 32'h68f02874;
    ram_cell[       4] = 32'h0;  // 32'he197d982;
    ram_cell[       5] = 32'h0;  // 32'h9928fa67;
    ram_cell[       6] = 32'h0;  // 32'hd7c0a01f;
    ram_cell[       7] = 32'h0;  // 32'h62fa5605;
    ram_cell[       8] = 32'h0;  // 32'h41c65a07;
    ram_cell[       9] = 32'h0;  // 32'h1b812f5d;
    ram_cell[      10] = 32'h0;  // 32'h07fcb0cb;
    ram_cell[      11] = 32'h0;  // 32'h79f07a8a;
    ram_cell[      12] = 32'h0;  // 32'h329ddb5e;
    ram_cell[      13] = 32'h0;  // 32'he202dd95;
    ram_cell[      14] = 32'h0;  // 32'hb0e41be8;
    ram_cell[      15] = 32'h0;  // 32'h1bdfe5bb;
    ram_cell[      16] = 32'h0;  // 32'hfae7186c;
    ram_cell[      17] = 32'h0;  // 32'h0972fbe5;
    ram_cell[      18] = 32'h0;  // 32'h26fcb26c;
    ram_cell[      19] = 32'h0;  // 32'ha0f48118;
    ram_cell[      20] = 32'h0;  // 32'h7ec3bb61;
    ram_cell[      21] = 32'h0;  // 32'hf90c709e;
    ram_cell[      22] = 32'h0;  // 32'hc1070330;
    ram_cell[      23] = 32'h0;  // 32'h98a926ff;
    ram_cell[      24] = 32'h0;  // 32'h50f9ace4;
    ram_cell[      25] = 32'h0;  // 32'ha9012651;
    ram_cell[      26] = 32'h0;  // 32'he1552907;
    ram_cell[      27] = 32'h0;  // 32'h683b05b0;
    ram_cell[      28] = 32'h0;  // 32'hf79d7ddb;
    ram_cell[      29] = 32'h0;  // 32'haadcbf56;
    ram_cell[      30] = 32'h0;  // 32'ha5462d94;
    ram_cell[      31] = 32'h0;  // 32'hc9b4c149;
    ram_cell[      32] = 32'h0;  // 32'h5b242abc;
    ram_cell[      33] = 32'h0;  // 32'hee0efd21;
    ram_cell[      34] = 32'h0;  // 32'h420eb9f1;
    ram_cell[      35] = 32'h0;  // 32'h73cf5ea3;
    ram_cell[      36] = 32'h0;  // 32'h7fcd4e99;
    ram_cell[      37] = 32'h0;  // 32'h507982e9;
    ram_cell[      38] = 32'h0;  // 32'hf2001510;
    ram_cell[      39] = 32'h0;  // 32'hf480a990;
    ram_cell[      40] = 32'h0;  // 32'ha9413b62;
    ram_cell[      41] = 32'h0;  // 32'h5bd939b6;
    ram_cell[      42] = 32'h0;  // 32'h01409a3c;
    ram_cell[      43] = 32'h0;  // 32'h22078c1f;
    ram_cell[      44] = 32'h0;  // 32'h30091e7e;
    ram_cell[      45] = 32'h0;  // 32'h825632f4;
    ram_cell[      46] = 32'h0;  // 32'he867ac9b;
    ram_cell[      47] = 32'h0;  // 32'h75c95a59;
    ram_cell[      48] = 32'h0;  // 32'heb4fd98c;
    ram_cell[      49] = 32'h0;  // 32'h6a6658f2;
    ram_cell[      50] = 32'h0;  // 32'he94d4a8b;
    ram_cell[      51] = 32'h0;  // 32'h79413027;
    ram_cell[      52] = 32'h0;  // 32'hddd3c7db;
    ram_cell[      53] = 32'h0;  // 32'he7818d37;
    ram_cell[      54] = 32'h0;  // 32'ha239e40b;
    ram_cell[      55] = 32'h0;  // 32'hd44a746e;
    ram_cell[      56] = 32'h0;  // 32'haf951834;
    ram_cell[      57] = 32'h0;  // 32'h1146b65b;
    ram_cell[      58] = 32'h0;  // 32'h4fd3085f;
    ram_cell[      59] = 32'h0;  // 32'hc804b838;
    ram_cell[      60] = 32'h0;  // 32'ha773834e;
    ram_cell[      61] = 32'h0;  // 32'h868111a7;
    ram_cell[      62] = 32'h0;  // 32'ha318f531;
    ram_cell[      63] = 32'h0;  // 32'h03483015;
    ram_cell[      64] = 32'h0;  // 32'h2fdbbad8;
    ram_cell[      65] = 32'h0;  // 32'h5b00c45e;
    ram_cell[      66] = 32'h0;  // 32'h4451bd99;
    ram_cell[      67] = 32'h0;  // 32'hca091efa;
    ram_cell[      68] = 32'h0;  // 32'h25a98b37;
    ram_cell[      69] = 32'h0;  // 32'hbee27df4;
    ram_cell[      70] = 32'h0;  // 32'h4aceeb34;
    ram_cell[      71] = 32'h0;  // 32'hd6062aaa;
    ram_cell[      72] = 32'h0;  // 32'hdff64303;
    ram_cell[      73] = 32'h0;  // 32'h3e51dd50;
    ram_cell[      74] = 32'h0;  // 32'h59ea79cf;
    ram_cell[      75] = 32'h0;  // 32'hf2489ec7;
    ram_cell[      76] = 32'h0;  // 32'hd79508e5;
    ram_cell[      77] = 32'h0;  // 32'h876d3151;
    ram_cell[      78] = 32'h0;  // 32'h08ce85a8;
    ram_cell[      79] = 32'h0;  // 32'h271b74b7;
    ram_cell[      80] = 32'h0;  // 32'h047ce3ac;
    ram_cell[      81] = 32'h0;  // 32'h970d3c55;
    ram_cell[      82] = 32'h0;  // 32'h7d909195;
    ram_cell[      83] = 32'h0;  // 32'h1d8acd6c;
    ram_cell[      84] = 32'h0;  // 32'h9c93eade;
    ram_cell[      85] = 32'h0;  // 32'h9398fea4;
    ram_cell[      86] = 32'h0;  // 32'hc852e9fb;
    ram_cell[      87] = 32'h0;  // 32'hf6c82001;
    ram_cell[      88] = 32'h0;  // 32'h2344d1dd;
    ram_cell[      89] = 32'h0;  // 32'h0c67857a;
    ram_cell[      90] = 32'h0;  // 32'h99fcaad5;
    ram_cell[      91] = 32'h0;  // 32'h8782d7a9;
    ram_cell[      92] = 32'h0;  // 32'h761e55d9;
    ram_cell[      93] = 32'h0;  // 32'he2e13597;
    ram_cell[      94] = 32'h0;  // 32'h1fb8c6bd;
    ram_cell[      95] = 32'h0;  // 32'h964d3df8;
    ram_cell[      96] = 32'h0;  // 32'hf53b10a9;
    ram_cell[      97] = 32'h0;  // 32'hd5f1d1e9;
    ram_cell[      98] = 32'h0;  // 32'h22ed277b;
    ram_cell[      99] = 32'h0;  // 32'h335b87de;
    ram_cell[     100] = 32'h0;  // 32'h74defff9;
    ram_cell[     101] = 32'h0;  // 32'hdacbbab0;
    ram_cell[     102] = 32'h0;  // 32'hfb0b9e8f;
    ram_cell[     103] = 32'h0;  // 32'h5ce7a697;
    ram_cell[     104] = 32'h0;  // 32'h64393860;
    ram_cell[     105] = 32'h0;  // 32'hcbabe1e4;
    ram_cell[     106] = 32'h0;  // 32'h2e1ef917;
    ram_cell[     107] = 32'h0;  // 32'h76a1e8e1;
    ram_cell[     108] = 32'h0;  // 32'hdf8fb853;
    ram_cell[     109] = 32'h0;  // 32'hfce528f2;
    ram_cell[     110] = 32'h0;  // 32'h7a844f03;
    ram_cell[     111] = 32'h0;  // 32'he44e2dab;
    ram_cell[     112] = 32'h0;  // 32'hc906c578;
    ram_cell[     113] = 32'h0;  // 32'h5fef0974;
    ram_cell[     114] = 32'h0;  // 32'hf12d9fb8;
    ram_cell[     115] = 32'h0;  // 32'h4d243983;
    ram_cell[     116] = 32'h0;  // 32'h62b6494e;
    ram_cell[     117] = 32'h0;  // 32'h2bef0b28;
    ram_cell[     118] = 32'h0;  // 32'hc7cfc8d3;
    ram_cell[     119] = 32'h0;  // 32'h803ae2da;
    ram_cell[     120] = 32'h0;  // 32'h91dc736a;
    ram_cell[     121] = 32'h0;  // 32'h351f1ae1;
    ram_cell[     122] = 32'h0;  // 32'h56b306e9;
    ram_cell[     123] = 32'h0;  // 32'h0e023ccd;
    ram_cell[     124] = 32'h0;  // 32'h0e8cd49e;
    ram_cell[     125] = 32'h0;  // 32'h7b806530;
    ram_cell[     126] = 32'h0;  // 32'h923d9646;
    ram_cell[     127] = 32'h0;  // 32'hd13d0240;
    ram_cell[     128] = 32'h0;  // 32'h118fa89c;
    ram_cell[     129] = 32'h0;  // 32'h60b0c933;
    ram_cell[     130] = 32'h0;  // 32'hb0446ab6;
    ram_cell[     131] = 32'h0;  // 32'h5235cd05;
    ram_cell[     132] = 32'h0;  // 32'hca51efa6;
    ram_cell[     133] = 32'h0;  // 32'h9a3a91c3;
    ram_cell[     134] = 32'h0;  // 32'h9c7fad0d;
    ram_cell[     135] = 32'h0;  // 32'h11a6c816;
    ram_cell[     136] = 32'h0;  // 32'hff8c3f32;
    ram_cell[     137] = 32'h0;  // 32'h0c90feb1;
    ram_cell[     138] = 32'h0;  // 32'h4e0a4a38;
    ram_cell[     139] = 32'h0;  // 32'h2dc3f1ed;
    ram_cell[     140] = 32'h0;  // 32'h8838dc0c;
    ram_cell[     141] = 32'h0;  // 32'he223da47;
    ram_cell[     142] = 32'h0;  // 32'h2e0353b1;
    ram_cell[     143] = 32'h0;  // 32'hd7aba25d;
    ram_cell[     144] = 32'h0;  // 32'hc86b2a4b;
    ram_cell[     145] = 32'h0;  // 32'h8215cd19;
    ram_cell[     146] = 32'h0;  // 32'h8f18281c;
    ram_cell[     147] = 32'h0;  // 32'h897ba662;
    ram_cell[     148] = 32'h0;  // 32'h477c347d;
    ram_cell[     149] = 32'h0;  // 32'h244745b2;
    ram_cell[     150] = 32'h0;  // 32'h8beabf19;
    ram_cell[     151] = 32'h0;  // 32'hc2f92d73;
    ram_cell[     152] = 32'h0;  // 32'hecfa1fe1;
    ram_cell[     153] = 32'h0;  // 32'hfee55d4a;
    ram_cell[     154] = 32'h0;  // 32'h40dfaedf;
    ram_cell[     155] = 32'h0;  // 32'hfab3e0b4;
    ram_cell[     156] = 32'h0;  // 32'h6344d432;
    ram_cell[     157] = 32'h0;  // 32'hc122b1c3;
    ram_cell[     158] = 32'h0;  // 32'h094ec522;
    ram_cell[     159] = 32'h0;  // 32'h6bf04b0e;
    ram_cell[     160] = 32'h0;  // 32'h8f7f4515;
    ram_cell[     161] = 32'h0;  // 32'h157e1e2a;
    ram_cell[     162] = 32'h0;  // 32'h59f934f1;
    ram_cell[     163] = 32'h0;  // 32'hbcafb3d9;
    ram_cell[     164] = 32'h0;  // 32'hb41a76e6;
    ram_cell[     165] = 32'h0;  // 32'h1d1be679;
    ram_cell[     166] = 32'h0;  // 32'h23d6a7e7;
    ram_cell[     167] = 32'h0;  // 32'he7244c44;
    ram_cell[     168] = 32'h0;  // 32'h2cd31f8a;
    ram_cell[     169] = 32'h0;  // 32'he33e3da4;
    ram_cell[     170] = 32'h0;  // 32'hfd055b0d;
    ram_cell[     171] = 32'h0;  // 32'hf08c1a3b;
    ram_cell[     172] = 32'h0;  // 32'hbd478de9;
    ram_cell[     173] = 32'h0;  // 32'hd4484841;
    ram_cell[     174] = 32'h0;  // 32'he300f934;
    ram_cell[     175] = 32'h0;  // 32'he7c53151;
    ram_cell[     176] = 32'h0;  // 32'h239820a3;
    ram_cell[     177] = 32'h0;  // 32'h6515396f;
    ram_cell[     178] = 32'h0;  // 32'had1712b2;
    ram_cell[     179] = 32'h0;  // 32'h9a6bfbe2;
    ram_cell[     180] = 32'h0;  // 32'h8c5f4c13;
    ram_cell[     181] = 32'h0;  // 32'h914ca497;
    ram_cell[     182] = 32'h0;  // 32'h49c76540;
    ram_cell[     183] = 32'h0;  // 32'hfe97a02a;
    ram_cell[     184] = 32'h0;  // 32'h1bc5d487;
    ram_cell[     185] = 32'h0;  // 32'h34dbbf6a;
    ram_cell[     186] = 32'h0;  // 32'h62b4c4a8;
    ram_cell[     187] = 32'h0;  // 32'h9d2008ee;
    ram_cell[     188] = 32'h0;  // 32'ha10d65e4;
    ram_cell[     189] = 32'h0;  // 32'hd64f5070;
    ram_cell[     190] = 32'h0;  // 32'hdf987e03;
    ram_cell[     191] = 32'h0;  // 32'h0d25c93b;
    ram_cell[     192] = 32'h0;  // 32'h60d3fdd3;
    ram_cell[     193] = 32'h0;  // 32'h35d1a5d2;
    ram_cell[     194] = 32'h0;  // 32'hb2f378a9;
    ram_cell[     195] = 32'h0;  // 32'h16daca16;
    ram_cell[     196] = 32'h0;  // 32'h36856fd2;
    ram_cell[     197] = 32'h0;  // 32'h384ab4ea;
    ram_cell[     198] = 32'h0;  // 32'h71bf4ce3;
    ram_cell[     199] = 32'h0;  // 32'h0877f8ce;
    ram_cell[     200] = 32'h0;  // 32'h30bf9860;
    ram_cell[     201] = 32'h0;  // 32'h3fb32cd8;
    ram_cell[     202] = 32'h0;  // 32'hedf36a09;
    ram_cell[     203] = 32'h0;  // 32'h2ed9b85d;
    ram_cell[     204] = 32'h0;  // 32'h539a513c;
    ram_cell[     205] = 32'h0;  // 32'h6ef47b0c;
    ram_cell[     206] = 32'h0;  // 32'hded949fc;
    ram_cell[     207] = 32'h0;  // 32'h4891a117;
    ram_cell[     208] = 32'h0;  // 32'h2655abe3;
    ram_cell[     209] = 32'h0;  // 32'h63ee326b;
    ram_cell[     210] = 32'h0;  // 32'h08aa0345;
    ram_cell[     211] = 32'h0;  // 32'h69cb48e0;
    ram_cell[     212] = 32'h0;  // 32'hd40a86b1;
    ram_cell[     213] = 32'h0;  // 32'hc3c07f79;
    ram_cell[     214] = 32'h0;  // 32'h7ec9c59f;
    ram_cell[     215] = 32'h0;  // 32'hd301abf0;
    ram_cell[     216] = 32'h0;  // 32'h3332e8b8;
    ram_cell[     217] = 32'h0;  // 32'h8e90a7e7;
    ram_cell[     218] = 32'h0;  // 32'hecde254e;
    ram_cell[     219] = 32'h0;  // 32'h3289794f;
    ram_cell[     220] = 32'h0;  // 32'ha5f025b0;
    ram_cell[     221] = 32'h0;  // 32'h43590ab5;
    ram_cell[     222] = 32'h0;  // 32'h6d118071;
    ram_cell[     223] = 32'h0;  // 32'h9fb47f68;
    ram_cell[     224] = 32'h0;  // 32'he9e3421f;
    ram_cell[     225] = 32'h0;  // 32'hd75605ff;
    ram_cell[     226] = 32'h0;  // 32'heeca00f9;
    ram_cell[     227] = 32'h0;  // 32'ha90bb137;
    ram_cell[     228] = 32'h0;  // 32'h56a6c480;
    ram_cell[     229] = 32'h0;  // 32'h8a9d2d9b;
    ram_cell[     230] = 32'h0;  // 32'h9072a501;
    ram_cell[     231] = 32'h0;  // 32'hbd578537;
    ram_cell[     232] = 32'h0;  // 32'h95525af6;
    ram_cell[     233] = 32'h0;  // 32'hf7dd0b45;
    ram_cell[     234] = 32'h0;  // 32'h88b06943;
    ram_cell[     235] = 32'h0;  // 32'h7e24facc;
    ram_cell[     236] = 32'h0;  // 32'h31394c20;
    ram_cell[     237] = 32'h0;  // 32'hf758a23d;
    ram_cell[     238] = 32'h0;  // 32'hd8a41bae;
    ram_cell[     239] = 32'h0;  // 32'h6f2bdcf8;
    ram_cell[     240] = 32'h0;  // 32'hbdc96eb1;
    ram_cell[     241] = 32'h0;  // 32'h57649298;
    ram_cell[     242] = 32'h0;  // 32'h6e8c8ba5;
    ram_cell[     243] = 32'h0;  // 32'hc6abe18a;
    ram_cell[     244] = 32'h0;  // 32'hc688ec36;
    ram_cell[     245] = 32'h0;  // 32'h26427e12;
    ram_cell[     246] = 32'h0;  // 32'h39fad76f;
    ram_cell[     247] = 32'h0;  // 32'hdde9e9de;
    ram_cell[     248] = 32'h0;  // 32'h9bc5de68;
    ram_cell[     249] = 32'h0;  // 32'h0566de1f;
    ram_cell[     250] = 32'h0;  // 32'hec8e067c;
    ram_cell[     251] = 32'h0;  // 32'h84857cf7;
    ram_cell[     252] = 32'h0;  // 32'hadef2d0b;
    ram_cell[     253] = 32'h0;  // 32'hf3178195;
    ram_cell[     254] = 32'h0;  // 32'hc3479240;
    ram_cell[     255] = 32'h0;  // 32'h2654abaf;
    // src matrix A
    ram_cell[     256] = 32'hbccde4ca;
    ram_cell[     257] = 32'h46fed4b9;
    ram_cell[     258] = 32'h6cdc03b7;
    ram_cell[     259] = 32'h62fb6370;
    ram_cell[     260] = 32'h42c6454c;
    ram_cell[     261] = 32'h971f004f;
    ram_cell[     262] = 32'he58aacb2;
    ram_cell[     263] = 32'h7badfe85;
    ram_cell[     264] = 32'h80408615;
    ram_cell[     265] = 32'h5b7c32f0;
    ram_cell[     266] = 32'hbf37743c;
    ram_cell[     267] = 32'h6bf9b3cc;
    ram_cell[     268] = 32'h1fdc9524;
    ram_cell[     269] = 32'h00651e74;
    ram_cell[     270] = 32'hc8f7f815;
    ram_cell[     271] = 32'hf5211de4;
    ram_cell[     272] = 32'h552d8977;
    ram_cell[     273] = 32'h040fac29;
    ram_cell[     274] = 32'ha73e0731;
    ram_cell[     275] = 32'h29b40822;
    ram_cell[     276] = 32'h370fffb1;
    ram_cell[     277] = 32'hc6c7b73b;
    ram_cell[     278] = 32'h1597467c;
    ram_cell[     279] = 32'h406a158c;
    ram_cell[     280] = 32'h0b3610b2;
    ram_cell[     281] = 32'h9e6977e1;
    ram_cell[     282] = 32'hae8cb1ea;
    ram_cell[     283] = 32'h5edb54b5;
    ram_cell[     284] = 32'hcc16f62e;
    ram_cell[     285] = 32'h90d7480d;
    ram_cell[     286] = 32'hbc0b1d9c;
    ram_cell[     287] = 32'h4b4677d9;
    ram_cell[     288] = 32'h171a03d6;
    ram_cell[     289] = 32'h2dad3ddf;
    ram_cell[     290] = 32'h93a55ebb;
    ram_cell[     291] = 32'h835d5dd5;
    ram_cell[     292] = 32'h41be2294;
    ram_cell[     293] = 32'h0661ede5;
    ram_cell[     294] = 32'h5df0f06d;
    ram_cell[     295] = 32'h2ed02d21;
    ram_cell[     296] = 32'h6e22b5b6;
    ram_cell[     297] = 32'h50bd4908;
    ram_cell[     298] = 32'h0948eb43;
    ram_cell[     299] = 32'h76af0502;
    ram_cell[     300] = 32'hbded2729;
    ram_cell[     301] = 32'h993ff92d;
    ram_cell[     302] = 32'h63028e01;
    ram_cell[     303] = 32'h0e630fb8;
    ram_cell[     304] = 32'hb371abc7;
    ram_cell[     305] = 32'hd1be6397;
    ram_cell[     306] = 32'h2b6dee79;
    ram_cell[     307] = 32'h4992505e;
    ram_cell[     308] = 32'hba5182bb;
    ram_cell[     309] = 32'hb319c630;
    ram_cell[     310] = 32'h2f37316a;
    ram_cell[     311] = 32'h17ff0f52;
    ram_cell[     312] = 32'h2814efbc;
    ram_cell[     313] = 32'hca93c702;
    ram_cell[     314] = 32'hffe432d1;
    ram_cell[     315] = 32'h03f0d0b2;
    ram_cell[     316] = 32'h2b2a7c77;
    ram_cell[     317] = 32'h235ae6d2;
    ram_cell[     318] = 32'h327b1d78;
    ram_cell[     319] = 32'h33c3a1a2;
    ram_cell[     320] = 32'h27bbadc9;
    ram_cell[     321] = 32'h544e4aa8;
    ram_cell[     322] = 32'he4b4a1a3;
    ram_cell[     323] = 32'h01dd258f;
    ram_cell[     324] = 32'hbc177725;
    ram_cell[     325] = 32'ha42e6b01;
    ram_cell[     326] = 32'h98a8d96c;
    ram_cell[     327] = 32'h1d11019f;
    ram_cell[     328] = 32'hf5d512b0;
    ram_cell[     329] = 32'hb15f92b3;
    ram_cell[     330] = 32'h95249981;
    ram_cell[     331] = 32'hf9b0d92c;
    ram_cell[     332] = 32'ha577103f;
    ram_cell[     333] = 32'h8facd16b;
    ram_cell[     334] = 32'h41aa6ffd;
    ram_cell[     335] = 32'h621ccd07;
    ram_cell[     336] = 32'h8579314a;
    ram_cell[     337] = 32'h59c51735;
    ram_cell[     338] = 32'hc8bfcdd2;
    ram_cell[     339] = 32'h91180f01;
    ram_cell[     340] = 32'hde300177;
    ram_cell[     341] = 32'hc403405b;
    ram_cell[     342] = 32'h88652f1b;
    ram_cell[     343] = 32'ha3bced2d;
    ram_cell[     344] = 32'h4ff02559;
    ram_cell[     345] = 32'h75653353;
    ram_cell[     346] = 32'hb063e26a;
    ram_cell[     347] = 32'h06506b3f;
    ram_cell[     348] = 32'he9130882;
    ram_cell[     349] = 32'h6c243fb1;
    ram_cell[     350] = 32'he711fdf3;
    ram_cell[     351] = 32'hdb084eab;
    ram_cell[     352] = 32'hdda58982;
    ram_cell[     353] = 32'h268f33b0;
    ram_cell[     354] = 32'h285972d4;
    ram_cell[     355] = 32'hb8a368bc;
    ram_cell[     356] = 32'hd8131145;
    ram_cell[     357] = 32'h8b3fc49c;
    ram_cell[     358] = 32'h39da5756;
    ram_cell[     359] = 32'hc0a4fc5b;
    ram_cell[     360] = 32'h675016af;
    ram_cell[     361] = 32'hee62213b;
    ram_cell[     362] = 32'h9452ab57;
    ram_cell[     363] = 32'h15b799c6;
    ram_cell[     364] = 32'h8adfbe3d;
    ram_cell[     365] = 32'h6698c810;
    ram_cell[     366] = 32'hbfc9f4a5;
    ram_cell[     367] = 32'h5da5cacd;
    ram_cell[     368] = 32'h1337f5c1;
    ram_cell[     369] = 32'h03d68b40;
    ram_cell[     370] = 32'h7ca79dae;
    ram_cell[     371] = 32'h2c482e3b;
    ram_cell[     372] = 32'h076f3f20;
    ram_cell[     373] = 32'ha5982e03;
    ram_cell[     374] = 32'h053bacd3;
    ram_cell[     375] = 32'h3799ebc1;
    ram_cell[     376] = 32'h50e3955d;
    ram_cell[     377] = 32'h450e8d08;
    ram_cell[     378] = 32'h5f0c67f1;
    ram_cell[     379] = 32'h478dcc1d;
    ram_cell[     380] = 32'h6db7a589;
    ram_cell[     381] = 32'hcf852738;
    ram_cell[     382] = 32'h3d954052;
    ram_cell[     383] = 32'h2111e710;
    ram_cell[     384] = 32'h3ad27e70;
    ram_cell[     385] = 32'h77d15836;
    ram_cell[     386] = 32'h04879f6a;
    ram_cell[     387] = 32'h6383c0c0;
    ram_cell[     388] = 32'h8402310f;
    ram_cell[     389] = 32'hdd4f2e57;
    ram_cell[     390] = 32'h02d3269a;
    ram_cell[     391] = 32'h5b5f975f;
    ram_cell[     392] = 32'hb364c03e;
    ram_cell[     393] = 32'hb3a4f488;
    ram_cell[     394] = 32'h999f5c0b;
    ram_cell[     395] = 32'h0d549b5a;
    ram_cell[     396] = 32'ha78abbe6;
    ram_cell[     397] = 32'h5f8a2ef9;
    ram_cell[     398] = 32'h65b0bb01;
    ram_cell[     399] = 32'h31b77936;
    ram_cell[     400] = 32'hc18ef873;
    ram_cell[     401] = 32'h7817ad6c;
    ram_cell[     402] = 32'h65009082;
    ram_cell[     403] = 32'h504d3449;
    ram_cell[     404] = 32'h4a8f05c2;
    ram_cell[     405] = 32'h01b17b1e;
    ram_cell[     406] = 32'h9606952d;
    ram_cell[     407] = 32'hdc36703d;
    ram_cell[     408] = 32'hd19c290b;
    ram_cell[     409] = 32'hb7d5207d;
    ram_cell[     410] = 32'h8b08c48d;
    ram_cell[     411] = 32'h02c34b80;
    ram_cell[     412] = 32'h45c6d087;
    ram_cell[     413] = 32'ha4d3ce37;
    ram_cell[     414] = 32'h6267dd8a;
    ram_cell[     415] = 32'h3c0142bc;
    ram_cell[     416] = 32'h2ca92ca4;
    ram_cell[     417] = 32'h65bb404f;
    ram_cell[     418] = 32'h97ec0b93;
    ram_cell[     419] = 32'h1d41c6bd;
    ram_cell[     420] = 32'h99cfef0d;
    ram_cell[     421] = 32'hb163f22f;
    ram_cell[     422] = 32'hcae544b3;
    ram_cell[     423] = 32'hbe69bc4a;
    ram_cell[     424] = 32'h8450b522;
    ram_cell[     425] = 32'h2c29bcce;
    ram_cell[     426] = 32'he3ed19f8;
    ram_cell[     427] = 32'h1b24e888;
    ram_cell[     428] = 32'h4552411d;
    ram_cell[     429] = 32'h96d70efa;
    ram_cell[     430] = 32'h0fcff269;
    ram_cell[     431] = 32'h74a4e8a5;
    ram_cell[     432] = 32'h226e5305;
    ram_cell[     433] = 32'he118a61a;
    ram_cell[     434] = 32'hb8893073;
    ram_cell[     435] = 32'heac83fb2;
    ram_cell[     436] = 32'had8d7590;
    ram_cell[     437] = 32'h587ca17a;
    ram_cell[     438] = 32'h6958900b;
    ram_cell[     439] = 32'hd8fdad9e;
    ram_cell[     440] = 32'h966e19d2;
    ram_cell[     441] = 32'h50d8e41c;
    ram_cell[     442] = 32'ha8ffb9c1;
    ram_cell[     443] = 32'h148e700b;
    ram_cell[     444] = 32'h4264a0f8;
    ram_cell[     445] = 32'hf3dd72db;
    ram_cell[     446] = 32'ha3384e6c;
    ram_cell[     447] = 32'h50e400c1;
    ram_cell[     448] = 32'h4b727853;
    ram_cell[     449] = 32'he788dd65;
    ram_cell[     450] = 32'h4a9193d8;
    ram_cell[     451] = 32'hf0675a89;
    ram_cell[     452] = 32'hce40ba1b;
    ram_cell[     453] = 32'hf2497124;
    ram_cell[     454] = 32'h6aeaa28a;
    ram_cell[     455] = 32'h53c03ecb;
    ram_cell[     456] = 32'hc116dbd5;
    ram_cell[     457] = 32'h20374821;
    ram_cell[     458] = 32'h9327e6ad;
    ram_cell[     459] = 32'h3443dd30;
    ram_cell[     460] = 32'hd562c73f;
    ram_cell[     461] = 32'h3adac98a;
    ram_cell[     462] = 32'hec614c89;
    ram_cell[     463] = 32'h740b3822;
    ram_cell[     464] = 32'hb36c3365;
    ram_cell[     465] = 32'h68dfbfbb;
    ram_cell[     466] = 32'h64f6c64f;
    ram_cell[     467] = 32'hb74e1389;
    ram_cell[     468] = 32'h10e74374;
    ram_cell[     469] = 32'he53f5a16;
    ram_cell[     470] = 32'ha32341de;
    ram_cell[     471] = 32'h04704783;
    ram_cell[     472] = 32'hc9acdb42;
    ram_cell[     473] = 32'hd64c7d4b;
    ram_cell[     474] = 32'hfde96d1e;
    ram_cell[     475] = 32'hd656f9e8;
    ram_cell[     476] = 32'hcde702fc;
    ram_cell[     477] = 32'hf97763d4;
    ram_cell[     478] = 32'h0b6c2963;
    ram_cell[     479] = 32'h132aaeaf;
    ram_cell[     480] = 32'hcc8f05c9;
    ram_cell[     481] = 32'hff788cd1;
    ram_cell[     482] = 32'hd8e24ac4;
    ram_cell[     483] = 32'h82187c7c;
    ram_cell[     484] = 32'hb50c7ae0;
    ram_cell[     485] = 32'h4bc4e43a;
    ram_cell[     486] = 32'h710f925f;
    ram_cell[     487] = 32'h278381aa;
    ram_cell[     488] = 32'hccd060a0;
    ram_cell[     489] = 32'hbbd930aa;
    ram_cell[     490] = 32'h359e3f78;
    ram_cell[     491] = 32'hef962d30;
    ram_cell[     492] = 32'hf4fd1a4b;
    ram_cell[     493] = 32'he8ac3533;
    ram_cell[     494] = 32'h9d55cf33;
    ram_cell[     495] = 32'h7410c98f;
    ram_cell[     496] = 32'h02c85f1b;
    ram_cell[     497] = 32'hde7dc724;
    ram_cell[     498] = 32'h312b6f7b;
    ram_cell[     499] = 32'hf99170f7;
    ram_cell[     500] = 32'h45c4f1b8;
    ram_cell[     501] = 32'h93702370;
    ram_cell[     502] = 32'haddeaad9;
    ram_cell[     503] = 32'h62f44495;
    ram_cell[     504] = 32'h49a0fe33;
    ram_cell[     505] = 32'h5049628a;
    ram_cell[     506] = 32'hf9a0d53a;
    ram_cell[     507] = 32'h0b3299df;
    ram_cell[     508] = 32'hfbe14397;
    ram_cell[     509] = 32'hccd97af3;
    ram_cell[     510] = 32'ha3a0998a;
    ram_cell[     511] = 32'h9c1ca68c;
    // src matrix B
    ram_cell[     512] = 32'h7c79527c;
    ram_cell[     513] = 32'h38573216;
    ram_cell[     514] = 32'h823a829e;
    ram_cell[     515] = 32'h18444b3b;
    ram_cell[     516] = 32'hb1643aec;
    ram_cell[     517] = 32'ha0497648;
    ram_cell[     518] = 32'h525ee633;
    ram_cell[     519] = 32'h0b32a9fe;
    ram_cell[     520] = 32'h68d73d7d;
    ram_cell[     521] = 32'hb38ae1fb;
    ram_cell[     522] = 32'hff1b143f;
    ram_cell[     523] = 32'hcf7e18c3;
    ram_cell[     524] = 32'hc6e94d32;
    ram_cell[     525] = 32'h60bc479e;
    ram_cell[     526] = 32'h17776e2e;
    ram_cell[     527] = 32'h835cbffc;
    ram_cell[     528] = 32'hbdd7b67a;
    ram_cell[     529] = 32'h2f8f8bb9;
    ram_cell[     530] = 32'hc2799da6;
    ram_cell[     531] = 32'h18b9a50f;
    ram_cell[     532] = 32'he91ebd8f;
    ram_cell[     533] = 32'ha543464b;
    ram_cell[     534] = 32'h4d43dd8d;
    ram_cell[     535] = 32'h39477433;
    ram_cell[     536] = 32'hc894676c;
    ram_cell[     537] = 32'h86384083;
    ram_cell[     538] = 32'h831ce9c5;
    ram_cell[     539] = 32'h1074dbd1;
    ram_cell[     540] = 32'hf705934b;
    ram_cell[     541] = 32'heba4d370;
    ram_cell[     542] = 32'h2bf7061e;
    ram_cell[     543] = 32'hea06912d;
    ram_cell[     544] = 32'hf776d660;
    ram_cell[     545] = 32'hb63ebff1;
    ram_cell[     546] = 32'h931279af;
    ram_cell[     547] = 32'h35d7ef40;
    ram_cell[     548] = 32'hfc392830;
    ram_cell[     549] = 32'h90c3725c;
    ram_cell[     550] = 32'h7f252fd4;
    ram_cell[     551] = 32'h541ac13c;
    ram_cell[     552] = 32'h53e5b396;
    ram_cell[     553] = 32'hb7b54daf;
    ram_cell[     554] = 32'h55de73fb;
    ram_cell[     555] = 32'he323c0ea;
    ram_cell[     556] = 32'h655633ca;
    ram_cell[     557] = 32'hfb075122;
    ram_cell[     558] = 32'h20fff5c5;
    ram_cell[     559] = 32'hf8683728;
    ram_cell[     560] = 32'h68f60437;
    ram_cell[     561] = 32'hd0a79203;
    ram_cell[     562] = 32'h57987b36;
    ram_cell[     563] = 32'h6adf1876;
    ram_cell[     564] = 32'he4a3953c;
    ram_cell[     565] = 32'h44660d04;
    ram_cell[     566] = 32'h481350f8;
    ram_cell[     567] = 32'ha98a62a7;
    ram_cell[     568] = 32'hd89211e8;
    ram_cell[     569] = 32'h42a3d80b;
    ram_cell[     570] = 32'ha567b646;
    ram_cell[     571] = 32'h5a3d0cbd;
    ram_cell[     572] = 32'h51f2caf5;
    ram_cell[     573] = 32'h9bc7d227;
    ram_cell[     574] = 32'h08d8a643;
    ram_cell[     575] = 32'he881b7df;
    ram_cell[     576] = 32'h138fa930;
    ram_cell[     577] = 32'h53ebd5bd;
    ram_cell[     578] = 32'h52ee8a0f;
    ram_cell[     579] = 32'hf4807de3;
    ram_cell[     580] = 32'h9928be97;
    ram_cell[     581] = 32'h26facc2e;
    ram_cell[     582] = 32'h323777f2;
    ram_cell[     583] = 32'h9e83dff8;
    ram_cell[     584] = 32'h7e4bb3b9;
    ram_cell[     585] = 32'h8e74fed6;
    ram_cell[     586] = 32'h1a1d89b2;
    ram_cell[     587] = 32'h686d7f74;
    ram_cell[     588] = 32'hccfc0f25;
    ram_cell[     589] = 32'hcedef876;
    ram_cell[     590] = 32'h4e77ae3b;
    ram_cell[     591] = 32'hdd1606ea;
    ram_cell[     592] = 32'h3e923eb2;
    ram_cell[     593] = 32'hf86c13f1;
    ram_cell[     594] = 32'hab84f218;
    ram_cell[     595] = 32'h43079003;
    ram_cell[     596] = 32'h749a4f81;
    ram_cell[     597] = 32'h18c3cbbd;
    ram_cell[     598] = 32'h432ab102;
    ram_cell[     599] = 32'h0fb9d9a0;
    ram_cell[     600] = 32'h806a22f6;
    ram_cell[     601] = 32'h231c5b3a;
    ram_cell[     602] = 32'h854e2fcb;
    ram_cell[     603] = 32'hdbac7a81;
    ram_cell[     604] = 32'h38fd03b5;
    ram_cell[     605] = 32'h29dca12c;
    ram_cell[     606] = 32'h46d02b18;
    ram_cell[     607] = 32'h5c2754bf;
    ram_cell[     608] = 32'h25f22c1d;
    ram_cell[     609] = 32'h15e6970c;
    ram_cell[     610] = 32'h8df114ac;
    ram_cell[     611] = 32'hb68f22c5;
    ram_cell[     612] = 32'h2267430b;
    ram_cell[     613] = 32'h65429555;
    ram_cell[     614] = 32'h55cf8864;
    ram_cell[     615] = 32'hba36133d;
    ram_cell[     616] = 32'h43e4d427;
    ram_cell[     617] = 32'h8d773501;
    ram_cell[     618] = 32'h21d4e24e;
    ram_cell[     619] = 32'hb6476473;
    ram_cell[     620] = 32'hc7104497;
    ram_cell[     621] = 32'h3c9bc61b;
    ram_cell[     622] = 32'h754d06c4;
    ram_cell[     623] = 32'h74cc05bb;
    ram_cell[     624] = 32'h802c5633;
    ram_cell[     625] = 32'hd6dd2c31;
    ram_cell[     626] = 32'h573e757d;
    ram_cell[     627] = 32'h26564551;
    ram_cell[     628] = 32'h65e23157;
    ram_cell[     629] = 32'hf152df6e;
    ram_cell[     630] = 32'he1f0d08b;
    ram_cell[     631] = 32'h82cc71ff;
    ram_cell[     632] = 32'hae4bafa2;
    ram_cell[     633] = 32'h2907e9cc;
    ram_cell[     634] = 32'h7478c788;
    ram_cell[     635] = 32'h5ac7b5a8;
    ram_cell[     636] = 32'h75077dd3;
    ram_cell[     637] = 32'h19b93881;
    ram_cell[     638] = 32'hff4651e9;
    ram_cell[     639] = 32'h97add7b6;
    ram_cell[     640] = 32'h1c058eaf;
    ram_cell[     641] = 32'h5925f357;
    ram_cell[     642] = 32'hd792f1c1;
    ram_cell[     643] = 32'h45610d57;
    ram_cell[     644] = 32'hbf5cf4b1;
    ram_cell[     645] = 32'h64335af2;
    ram_cell[     646] = 32'h22c27c4b;
    ram_cell[     647] = 32'h5ca26d38;
    ram_cell[     648] = 32'hbfe06a5e;
    ram_cell[     649] = 32'he3ea7471;
    ram_cell[     650] = 32'hffda0dc4;
    ram_cell[     651] = 32'h73e173f9;
    ram_cell[     652] = 32'hb6b0b7ea;
    ram_cell[     653] = 32'h45a39797;
    ram_cell[     654] = 32'hdf947b4a;
    ram_cell[     655] = 32'h1346af55;
    ram_cell[     656] = 32'h7f4ab182;
    ram_cell[     657] = 32'he74a78c2;
    ram_cell[     658] = 32'h2c1af989;
    ram_cell[     659] = 32'ha5e8bdc3;
    ram_cell[     660] = 32'h03ae8443;
    ram_cell[     661] = 32'h28a4ee96;
    ram_cell[     662] = 32'h04597bee;
    ram_cell[     663] = 32'h3662f441;
    ram_cell[     664] = 32'he2b77e3f;
    ram_cell[     665] = 32'h1d8b8fb8;
    ram_cell[     666] = 32'h214965b7;
    ram_cell[     667] = 32'h30e67a3c;
    ram_cell[     668] = 32'h8f4565d3;
    ram_cell[     669] = 32'h29f79757;
    ram_cell[     670] = 32'h03b2db14;
    ram_cell[     671] = 32'h6ec707ae;
    ram_cell[     672] = 32'h80001cc6;
    ram_cell[     673] = 32'hd30c3b41;
    ram_cell[     674] = 32'h1de77038;
    ram_cell[     675] = 32'h1106c3b1;
    ram_cell[     676] = 32'h68dcd233;
    ram_cell[     677] = 32'h8d5e1d72;
    ram_cell[     678] = 32'h1e0a79a9;
    ram_cell[     679] = 32'hbdeae96a;
    ram_cell[     680] = 32'h764ac524;
    ram_cell[     681] = 32'h4e0d2933;
    ram_cell[     682] = 32'he83f01a2;
    ram_cell[     683] = 32'h5a3cca6b;
    ram_cell[     684] = 32'h1e28711a;
    ram_cell[     685] = 32'h230f1720;
    ram_cell[     686] = 32'hd0aebca6;
    ram_cell[     687] = 32'hc9a9476b;
    ram_cell[     688] = 32'h7699c65e;
    ram_cell[     689] = 32'hc976a283;
    ram_cell[     690] = 32'h7a9dc585;
    ram_cell[     691] = 32'h908d8cae;
    ram_cell[     692] = 32'ha0ba9eed;
    ram_cell[     693] = 32'h1a6e194a;
    ram_cell[     694] = 32'h3fdad771;
    ram_cell[     695] = 32'hfc19e010;
    ram_cell[     696] = 32'h28a637a0;
    ram_cell[     697] = 32'h51b5e421;
    ram_cell[     698] = 32'h0755b7a3;
    ram_cell[     699] = 32'hd63b35e2;
    ram_cell[     700] = 32'hb9ba39a6;
    ram_cell[     701] = 32'h913162d9;
    ram_cell[     702] = 32'he8e73837;
    ram_cell[     703] = 32'h06a2e908;
    ram_cell[     704] = 32'hf984c186;
    ram_cell[     705] = 32'he2ee0544;
    ram_cell[     706] = 32'hcffe88d9;
    ram_cell[     707] = 32'hea029a7b;
    ram_cell[     708] = 32'h7a41c6f6;
    ram_cell[     709] = 32'he2abe946;
    ram_cell[     710] = 32'hefa4794a;
    ram_cell[     711] = 32'h2526fc3b;
    ram_cell[     712] = 32'h1a46750c;
    ram_cell[     713] = 32'h24b8907d;
    ram_cell[     714] = 32'he154cc44;
    ram_cell[     715] = 32'ha63ac651;
    ram_cell[     716] = 32'h4f717798;
    ram_cell[     717] = 32'h67dcb949;
    ram_cell[     718] = 32'h0f15b615;
    ram_cell[     719] = 32'h2090b251;
    ram_cell[     720] = 32'he35804c9;
    ram_cell[     721] = 32'heda4cd0d;
    ram_cell[     722] = 32'hd98a69f6;
    ram_cell[     723] = 32'he0393055;
    ram_cell[     724] = 32'h56111e42;
    ram_cell[     725] = 32'h3037ad45;
    ram_cell[     726] = 32'h5a53be9b;
    ram_cell[     727] = 32'h0cd072ba;
    ram_cell[     728] = 32'h9201cb4a;
    ram_cell[     729] = 32'h87d5dd84;
    ram_cell[     730] = 32'h00952327;
    ram_cell[     731] = 32'hd21bc190;
    ram_cell[     732] = 32'h8a9e356e;
    ram_cell[     733] = 32'h36be0815;
    ram_cell[     734] = 32'h3c55b7c1;
    ram_cell[     735] = 32'h199f3805;
    ram_cell[     736] = 32'h65b6fd00;
    ram_cell[     737] = 32'hc2e75528;
    ram_cell[     738] = 32'hee5318f8;
    ram_cell[     739] = 32'hd1b412ac;
    ram_cell[     740] = 32'h7f2ae33a;
    ram_cell[     741] = 32'h8961c797;
    ram_cell[     742] = 32'h248c9238;
    ram_cell[     743] = 32'h0b066699;
    ram_cell[     744] = 32'hb8ccdd03;
    ram_cell[     745] = 32'h9e4af888;
    ram_cell[     746] = 32'h0859f4aa;
    ram_cell[     747] = 32'hb3fb6433;
    ram_cell[     748] = 32'hfa19bc3f;
    ram_cell[     749] = 32'h4a46191d;
    ram_cell[     750] = 32'h92091518;
    ram_cell[     751] = 32'h9aa3946c;
    ram_cell[     752] = 32'hdafc1a0d;
    ram_cell[     753] = 32'h9bb66dff;
    ram_cell[     754] = 32'h79aff052;
    ram_cell[     755] = 32'heafb5124;
    ram_cell[     756] = 32'h687e6516;
    ram_cell[     757] = 32'ha28d737b;
    ram_cell[     758] = 32'hd06d2c44;
    ram_cell[     759] = 32'h0d0e6ce9;
    ram_cell[     760] = 32'h6574778f;
    ram_cell[     761] = 32'hd4cb929b;
    ram_cell[     762] = 32'h9fea301e;
    ram_cell[     763] = 32'h8d98c03f;
    ram_cell[     764] = 32'h93ba337b;
    ram_cell[     765] = 32'h1edf8a41;
    ram_cell[     766] = 32'h46de447c;
    ram_cell[     767] = 32'h6d4d64e8;
end

endmodule
